
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package prog_mem_content is

-- content of pe_0 ----------------------------------------------------------------------------------
constant pe_0_00 : BIT_VECTOR := X"033C94222AF38FC23C40FFFFF8F412492595C5550AEF128010C84E3579BDF135";
constant pe_0_01 : BIT_VECTOR := X"077870EBC9F960558E9D4489ACC80D8D85C8E0A19F9811A081F8F068DC8002AE";
constant pe_0_02 : BIT_VECTOR := X"8FFFFFFFFFFF33C3C1B0EE8E05BC9F950CC8C805C9B0D8C91A0D6C9F9A8C9F95";
constant pe_0_03 : BIT_VECTOR := X"7D10ED85F1B0FFDBEEA8F01F08DE8AD889D10ED87F1D0FFDBEEA8101F08DE8AD";
constant pe_0_04 : BIT_VECTOR := X"07F001242FF0010FF1F8010FF108EC1C1BA03EF981EA1E01D120F7F80DFFFFF8";
constant pe_0_05 : BIT_VECTOR := X"0FF7C179FB7C979FB6C269FB6CA69FB5C359FB5CB59FB4C449FB4CC49FB00C01";
constant pe_0_06 : BIT_VECTOR := X"0E04E00E0CFFDAEA51EE197969594939291909796959493929190080FC23B911";
constant pe_0_07 : BIT_VECTOR := X"C898808C08F08D08608B09D8A3C03C07C03E066E02E0C06E05C05C01C05E04E0";
constant pe_0_08 : BIT_VECTOR := X"87E8D765B445E4E74C4AB80F9E433A80F23A8E10F6AC205315732279B7F79B10";
constant pe_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6020C0C5923BD29";
constant pe_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_1 ----------------------------------------------------------------------------------
constant pe_1_00 : BIT_VECTOR := X"B1FFF333394F942AFF24C0ECAFBFEA0DA0F8003B4EDC10010DCCCDFFFFFFF002";
constant pe_1_01 : BIT_VECTOR := X"411A366FE118F111CC6E11CEEECDCC44444555E477BE11E445A0044556AABADB";
constant pe_1_02 : BIT_VECTOR := X"DD1FDACE0CFFF23FF2F4116344F518FF411A3EEF1D2CCFDDDFCCFD77BE6755AF";
constant pe_1_03 : BIT_VECTOR := X"F8088FF08801E8F1880018F88881108D138088FF48841E8F1880068F88881108";
constant pe_1_04 : BIT_VECTOR := X"28F0E898EFF80E28F78F0E28F88F0002E888CC648DC80DEE01F8810FECCDF1D1";
constant pe_1_05 : BIT_VECTOR := X"8D188A98BD88A98BD88A98BD88A98BD88A98BD88A98BD88A98BD88A98BDB8F0E";
constant pe_1_06 : BIT_VECTOR := X"8BB8BB8BBF1D16C126CC188888888888888888888888888888888E8992AFF288";
constant pe_1_07 : BIT_VECTOR := X"B888890890890890890890EF889AA9AA9AABB82BB2BB8AABB89AA9AA9AABB8BB";
constant pe_1_08 : BIT_VECTOR := X"288915FB87B2AF43EA230B941741FD34903A5BB02D52B8023EF97A4CA667F389";
constant pe_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF32036266677B248";
constant pe_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_2 ----------------------------------------------------------------------------------
constant pe_2_00 : BIT_VECTOR := X"07F1F77751D43F1FF1F033222417770770F1011103F54CE20333333333333440";
constant pe_2_01 : BIT_VECTOR := X"176E63510FF11176EE1576F11E11FDFF3711F010FF11761F191FF371F1FFF51F";
constant pe_2_02 : BIT_VECTOR := X"0332200011E5471F1F1176F63711F111176E63F11F63711EC03711FF1111FF11";
constant pe_2_03 : BIT_VECTOR := X"1D7756E2D7274547557F2F657755F5D472D7752E2D7270503553F2F657355F1D";
constant pe_2_04 : BIT_VECTOR := X"001000426AF107003101070031F1DF20C44101D03115012726010AE477300117";
constant pe_2_05 : BIT_VECTOR := X"13371957F131917F171957F131917F171957F131917F171957F131917F111107";
constant pe_2_06 : BIT_VECTOR := X"7F03F03F0111F010FF11075757575757575757171717171717171630F1FF1F01";
constant pe_2_07 : BIT_VECTOR := X"1F7F305C05705705605504E4031F11F11F5F073F03F01F1F071F51F51F1F07F0";
constant pe_2_08 : BIT_VECTOR := X"F941E9E6AF6E8A9D92CAB48C3D7C215F8F5BF9BD430A52A351C60F0D6B5BB200";
constant pe_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF04047C9F956F8D";
constant pe_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_3 ----------------------------------------------------------------------------------
constant pe_3_00 : BIT_VECTOR := X"E91019229029F590102E999999D0F1CF1929C999EEBE23001CCCCCCCCCCCCCCC";
constant pe_3_01 : BIT_VECTOR := X"8990982091400899000299000298520582984E05140099058000582849077904";
constant pe_3_02 : BIT_VECTOR := X"8999999999C19291050899098209100089909820919820911E82091400891400";
constant pe_3_03 : BIT_VECTOR := X"D222282D22D282882282D222282228282D222282D22D282882282D2222822282";
constant pe_3_04 : BIT_VECTOR := X"4EEC45EF10E80F4EED700F4EED7000EC2EEED05C2D0990EF99EEEBB99B999992";
constant pe_3_05 : BIT_VECTOR := X"999895824089582408958240895824089582408958240895824089582400E00F";
constant pe_3_06 : BIT_VECTOR := X"84E84E84E099DE03D200E28282828282828282828282828282828EFE590102E1";
constant pe_3_07 : BIT_VECTOR := X"00202E9EE9EE9EE9EE9EE95F389589589584E884E84E9584E89589589584E84E";
constant pe_3_08 : BIT_VECTOR := X"DE919B0681C20EA67650D18D731ED2F8A78FC35E8BA17E9C1FC2CAF772C7C0EE";
constant pe_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF40367676741060";
constant pe_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_0 ----------------------------------------------------------------------------------
constant po_0_00 : BIT_VECTOR := X"0CF20890020DF003B20BFFFFFF01B3DE3D8F575570D4F02B00EA621468ACE024";
constant po_0_01 : BIT_VECTOR := X"6AC9F980668A0E8C91580C948D33E09F9B22A081F8E85C8E0A29F957A09AA21C";
constant po_0_02 : BIT_VECTOR := X"9CFFF8FFFFF8A08F2F056C9F980DD8D01AC9F910BB8960AA8F9B099878788880";
constant po_0_03 : BIT_VECTOR := X"EEE8E01F0CDE8EDC88D10E986F1C0BF9FEEE8001F0CDE8EDC8AD10E988F1E0BF";
constant po_0_04 : BIT_VECTOR := X"011010FF10FC8001250080012500FD081A9581FE9211D120A1E014DEFEF8FFFF";
constant po_0_05 : BIT_VECTOR := X"BCF89FB3C539FB3CD39FB2C629FB2CE29FB1C719FB1CF19FB0C809FB0C018090";
constant po_0_06 : BIT_VECTOR := X"4C00C04C008F0E80FEA28FFEEDDCCBBAA9988FFEEDDCCBBAA99880B0103A204E";
constant po_0_07 : BIT_VECTOR := X"088B48608F08708D08F08FFC187E03E07E0C072C06C02E0C021E05E01E0C01C0";
constant po_0_08 : BIT_VECTOR := X"CEB916180B8CA5CD71290E62044FD0C210530AA0392B9B7841467CDAAE02380C";
constant po_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF08D0FF8E0E101F";
constant po_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_1 ----------------------------------------------------------------------------------
constant po_1_00 : BIT_VECTOR := X"AADEDEF2325FF42BDE30D1FDBF03EB1FB0EE902A1FCD180380CCCCCFFFFFF000";
constant po_1_01 : BIT_VECTOR := X"4F6B5FF6110011FEDDEEEDD2EE11DD55AE11E445A66444555E411844E4BBBB17";
constant po_1_02 : BIT_VECTOR := X"FEC0E0BDF1D0F221E344F57BFF4110344F1B5FE011CEFC11CC6FC11666611444";
constant po_1_03 : BIT_VECTOR := X"8800F8F88881108D118088FF28821E8F1880048F88881108D158088FF68861E8";
constant po_1_04 : BIT_VECTOR := X"8F20E9E8F2E8F08F2898108F28981111F888147B080E05F880DE81CD0DD0E0C1";
constant po_1_05 : BIT_VECTOR := X"3AC08BD88A98BD88A98BD88A98BD88A98BD88A98BD88A98BD88A98BD88A169A0";
constant po_1_06 : BIT_VECTOR := X"A8AA8AA8AA0C8C0B1C11089898989898989898989898989898989FE902BDE360";
constant po_1_07 : BIT_VECTOR := X"8009208908908908908908FF909BB9BB9BB8AA92AA2AABB9AA9BB9BB9BB8AA8A";
constant po_1_08 : BIT_VECTOR := X"8C96E86474E1B668E9C4ED4266C5C1B95544D46252510E010733B9AFCF3F6084";
constant po_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80836666766B4B";
constant po_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_2 ----------------------------------------------------------------------------------
constant po_2_00 : BIT_VECTOR := X"F11F0F1FF500413F1F0033222F07472172F11D1100F0E0B01033333333333444";
constant po_2_01 : BIT_VECTOR := X"711E111176FF3510EC0310F62676F0FF11761F191FF3711F010FF17F1DF77571";
constant po_2_02 : BIT_VECTOR := X"0133250001100316FF3711F111176F63711E117176F11176EE11176FF3776FF3";
constant po_2_03 : BIT_VECTOR := X"557F1F657755F5D472D7756E2D7274543553F2F657355F1D072D7752E2D72705";
constant po_2_04 : BIT_VECTOR := X"00A0700341A910004B01A0004B01DF0AC33BA6F1436726015011BAFF67350117";
constant po_2_05 : BIT_VECTOR := X"21357F171957F131917F171957F131917F171957F131917F171957F131A4F1F0";
constant po_2_06 : BIT_VECTOR := X"51F51F11F1510103F1E007575757575757575313131313131313101103F1F000";
constant po_2_07 : BIT_VECTOR := X"6551450056050056054053F1553F07F07F01F571F51F5F01F17F03F03F01F11F";
constant po_2_08 : BIT_VECTOR := X"15E98153EDD68A6585362EEA1D77CF6D3C9DFCBC13BE3726785FD449271BC53C";
constant po_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB0102C5B435496";
constant po_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_3 ----------------------------------------------------------------------------------
constant po_3_00 : BIT_VECTOR := X"5900800779EC238100EC99999CCF309009209F99CEBEB03006CCCCCCCCCCCCCC";
constant po_3_01 : BIT_VECTOR := X"209100089905820911E8891982994E140099058000582984E051402205122999";
constant po_3_02 : BIT_VECTOR := X"80999999999FE889048209100089909820910028990008990000899058299058";
constant po_3_03 : BIT_VECTOR := X"2282D222282228282D222282D22D282882282D222282228282D222282D22D282";
constant po_3_04 : BIT_VECTOR := X"45E0F4EE0E1B0C45EBE8BC45EBE811EB2AABB940FB9F99EE990EBBBBBB999998";
constant po_3_05 : BIT_VECTOR := X"00992408958240895824089582408958240895824089582408958240895298CC";
constant po_3_06 : BIT_VECTOR := X"895895895899E0DF50DDC88888888888888888888888888888888E03C8100ECC";
constant po_3_07 : BIT_VECTOR := X"E99EF9EE9EE9EE9EE9EE9E400984E84E84E95889589584E95884E84E84E95895";
constant po_3_08 : BIT_VECTOR := X"A51DFC303BDA775DC9D035E285A90FB9A3F4E4CFDE368219CDA3FAD58D06799D";
constant po_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1103726476659E";
constant po_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

end prog_mem_content;



library IEEE;
use IEEE.STD_LOGIC_1164.all;

package prog_mem_content is

-- content of pe_0 ----------------------------------------------------------------------------------
constant pe_0_00 : BIT_VECTOR := X"002AE033C94222AF38FC23C40FFFFF89412492595C55506EF1270168ACE0246B";
constant pe_0_01 : BIT_VECTOR := X"C9F95077870EBC9F960558E9D4489ACC80D8D85C8E0A19F9811A081F8F068DC8";
constant pe_0_02 : BIT_VECTOR := X"DE8AD8FFFFFFFFFFF33C3C1B0EE8E05BC9F950CC8C805C9B0D8C91A0D6C9F9A8";
constant pe_0_03 : BIT_VECTOR := X"FFFF84D10ED82F180FFDBEEA8C01F08DE8AD886D10ED84F1A0FFDBEEA8E01F08";
constant pe_0_04 : BIT_VECTOR := X"110FF7C179FB7C979FB6C269FB6CA69FB5C359FB5CB59FB4C449FB4CC49FB00C";
constant pe_0_05 : BIT_VECTOR := X"E00E04E00E0CFFDAEA51EE197969594939291909796959493929190080FC23B9";
constant pe_0_06 : BIT_VECTOR := X"8B4800117EE88880E564347E00F3C03C07C03E066E02E0C06E05C05C01C05E04";
constant pe_0_07 : BIT_VECTOR := X"B916180B8CA5CD71290E62044FD0C210530AA0392B9B7841467CDAAE02380F08";
constant pe_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF08D01FCE";
constant pe_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_1 ----------------------------------------------------------------------------------
constant pe_1_00 : BIT_VECTOR := X"ABADBB1FFF333394F942AFF24C0ECAF0FEA0DA0F8003B4EDC100107777788881";
constant pe_1_01 : BIT_VECTOR := X"755AF411A366FE118F111CC6E11CEEECDCC44444555E477BE11E445A0044556A";
constant pe_1_02 : BIT_VECTOR := X"81108DD1FDACE0CFFF23FF2F4116344F518FF411A3EEF1D2CCFDDDFCCFD77BE6";
constant pe_1_03 : BIT_VECTOR := X"DF1D188088FF98891E8F18800A8F88881108D1C8088FFD88D1E8F18800E8F888";
constant pe_1_04 : BIT_VECTOR := X"888D188A98BD88A98BD88A98BD88A98BD88A98BD88A98BD88A98BD88A98BDB8F";
constant pe_1_05 : BIT_VECTOR := X"BB8BB8BB8BBF1D16C126CC188888888888888888888888888888888E8992AFF2";
constant pe_1_06 : BIT_VECTOR := X"092E09280C680882C888888D00C89AA9AA9AABB82BB2BB8AABB89AA9AA9AABB8";
constant pe_1_07 : BIT_VECTOR := X"96E86474E1B668E9C4ED4266C5C1B95544D46252510E010733B9AFCF3F608B80";
constant pe_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF808B4B8C";
constant pe_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_2 ----------------------------------------------------------------------------------
constant pe_2_00 : BIT_VECTOR := X"FF51F07F1F77751D43F1FF1F033222437770770F1011102F54C4203333333330";
constant pe_2_01 : BIT_VECTOR := X"1FF11176E63510FF11176EE1576F11E11FDFF3711F010FF11761F191FF371F1F";
constant pe_2_02 : BIT_VECTOR := X"55F1D0332200011E5471F1F1176F63711F111176E63F11F63711EC03711FF111";
constant pe_2_03 : BIT_VECTOR := X"001171D7756E1D7174547557F1F657755F5D471D7752E1D7170503553F1F6573";
constant pe_2_04 : BIT_VECTOR := X"0113371957F131917F171957F131917F171957F131917F171957F131917F1111";
constant pe_2_05 : BIT_VECTOR := X"F07F03F03F0111F010FF11075757575757575757171717171717171630F1FF1F";
constant pe_2_06 : BIT_VECTOR := X"514F000EF1FB083010000BB700331F11F11F5F073F03F01F1F071F51F51F1F07";
constant pe_2_07 : BIT_VECTOR := X"E98153EDD68A6585362EEA1D77CF6D3C9DFCBC13BE3726785FD449271BC53C65";
constant pe_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB0149615";
constant pe_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_3 ----------------------------------------------------------------------------------
constant pe_3_00 : BIT_VECTOR := X"77904E91019229029F590102E999999D0F1CF1929C999EEBE21101CCCCCCCCCC";
constant pe_3_01 : BIT_VECTOR := X"914008990982091400899000299000298520582984E051400990580005828490";
constant pe_3_02 : BIT_VECTOR := X"222828999999999C19291050899098209100089909820919820911E820914008";
constant pe_3_03 : BIT_VECTOR := X"99992D222282D22D282882282D222282228282D222282D22D282882282D22228";
constant pe_3_04 : BIT_VECTOR := X"E1999895824089582408958240895824089582408958240895824089582400E0";
constant pe_3_05 : BIT_VECTOR := X"4E84E84E84E099DE03D200E28282828282828282828282828282828EFE590102";
constant pe_3_06 : BIT_VECTOR := X"9EFCC45ED05BCE2D0EEEEBBBDD989589589584E884E84E9584E89589589584E8";
constant pe_3_07 : BIT_VECTOR := X"1DFC303BDA775DC9D035E285A90FB9A3F4E4CFDE368219CDA3FAD58D06799DE9";
constant pe_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF11059EA5";
constant pe_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_0 ----------------------------------------------------------------------------------
constant po_0_00 : BIT_VECTOR := X"AA21C0CF20890020DF003B20BFFFFFF0173DE3D8F575570D4F02B0079BDF1357";
constant po_0_01 : BIT_VECTOR := X"888806AC9F980668A0E8C91580C948D33E09F9B22A081F8E85C8E0A29F957A09";
constant po_0_02 : BIT_VECTOR := X"1B0BF9CFFF8FFFFF8A08F2F056C9F980DD8D01AC9F910BB8960AA8F9B0998787";
constant po_0_03 : BIT_VECTOR := X"8FFFFEEE8B01F0CDE8EDC85D10E983F190BF9FEEE8D01F0CDE8EDC87D10E985F";
constant po_0_04 : BIT_VECTOR := X"4EBCF89FB3C539FB3CD39FB2C629FB2CE29FB1C719FB1CF19FB0C809FB0C0180";
constant po_0_05 : BIT_VECTOR := X"C04C00C04C008F0E80FE428FFEEDDCCBBAA9988FFEEDDCCBBAA99880B0103A20";
constant po_0_06 : BIT_VECTOR := X"89880104F3FEF89519EDCB0FD0F87E03E07E0C072C06C02E0C021E05E01E0C01";
constant po_0_07 : BIT_VECTOR := X"7E8D765B445E4E74C4AB80F9E433A80F23A8E10F6AC205315732279B7F76B10C";
constant po_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF602BD298";
constant po_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_1 ----------------------------------------------------------------------------------
constant po_1_00 : BIT_VECTOR := X"BBB17AADEDEF2325FF42BDE30D1FDBF03EB1FB0EE902A1FCD180180777778888";
constant po_1_01 : BIT_VECTOR := X"114444F6B5FF6110011FEDDEEEDD2EE11DD55AE11E445A66444555E411844E4B";
constant po_1_02 : BIT_VECTOR := X"8F1E8FEC0E0BDF1D0F221E344F57BFF4110344F1B5FE011CEFC11CC6FC116666";
constant po_1_03 : BIT_VECTOR := X"0E0C1880088F88881108D1A8088FFB88B1E8F18800C8F88881108D1E8088FFF8";
constant po_1_04 : BIT_VECTOR := X"601AC08BD88A98BD88A98BD88A98BD88A98BD88A98BD88A98BD88A98BD88A169";
constant po_1_05 : BIT_VECTOR := X"8AA8AA8AA8AA0C8C0B1C91089898989898989898989898989898989FE902BDE3";
constant po_1_06 : BIT_VECTOR := X"88880E89207B881808888188C0D09BB9BB9BB8AA92AA2AABB9AA9BB9BB9BB8AA";
constant po_1_07 : BIT_VECTOR := X"88915FB87B2AF43EA230B941741FD34903A5BB02D52B8023EF97A4CA6677189B";
constant po_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF320B2482";
constant po_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_2 ----------------------------------------------------------------------------------
constant po_2_00 : BIT_VECTOR := X"77571F11F0F1FF500413F1F0033222F07372172F11D1100F0E0B010333333333";
constant po_2_01 : BIT_VECTOR := X"76FF3711E111176FF3510EC0310F62676F0FF11761F191FF3711F010FF17F1FF";
constant po_2_02 : BIT_VECTOR := X"717050133250001100316FF3711F111176F63711E117176F11176EE11176FF37";
constant po_2_03 : BIT_VECTOR := X"50117557F1F657755F5D471D7756E1D7174543553F1F657355F1D071D7752E1D";
constant po_2_04 : BIT_VECTOR := X"0021357F171957F131917F171957F131917F171957F131917F171957F131A4F1";
constant po_2_05 : BIT_VECTOR := X"1F51F51F11F1510103F1E007575757575757575313131313131313101103F1F0";
constant po_2_06 : BIT_VECTOR := X"F7F30700F6F17B03633332FF70353F07F07F01F571F51F5F01F17F03F03F01F1";
constant po_2_07 : BIT_VECTOR := X"941E9E6AF6E8A9D92CAB48C3D7C215F8F5BF9BD430A52A351C60F0D6B5BC2001";
constant po_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF046F8DF";
constant po_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_3 ----------------------------------------------------------------------------------
constant po_3_00 : BIT_VECTOR := X"229995900800779EC238100EC99999CCF309009209F99CEBEB01006CCCCCCCCC";
constant po_3_01 : BIT_VECTOR := X"99058209100089905820911E8891982994E140099058000582984E0514022051";
constant po_3_02 : BIT_VECTOR := X"2D28280999999999FE8890482091000899098209100289900089900008990582";
constant po_3_03 : BIT_VECTOR := X"999982282D222282228282D222282D22D282882282D222282228282D222282D2";
constant po_3_04 : BIT_VECTOR := X"CC00992408958240895824089582408958240895824089582408958240895298";
constant po_3_05 : BIT_VECTOR := X"95895895895899E0DF50DDC88888888888888888888888888888888E03C8100E";
constant po_3_06 : BIT_VECTOR := X"02020F4EE940EBFB988888EEBD9984E84E84E95889589584E95884E84E84E958";
constant po_3_07 : BIT_VECTOR := X"E919B0681C20EA67650D18D731ED2F8A78FC35E8BA17E9C1FC2CAF772C7C0EE0";
constant po_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF401060D";
constant po_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

end prog_mem_content;



library IEEE;
use IEEE.STD_LOGIC_1164.all;

package prog_mem_content is

-- content of pe_0 ----------------------------------------------------------------------------------
constant pe_0_00 : BIT_VECTOR := X"89049A89DFA409ADEFEFFFFFFFFF8A412492595C5550AEF101D95FACE02468AF";
constant pe_0_01 : BIT_VECTOR := X"EF71A99E97F333928581FF7380C06E01E31A688913210D0309001E65127949FF";
constant pe_0_02 : BIT_VECTOR := X"199C2F031F10A19E9019C318794912126FF7110690BF0E4F0320EF7FE64F0320";
constant pe_0_03 : BIT_VECTOR := X"8608D0060F64589104EB435E9B8936F58FEF700F7207220066A94D8519681510";
constant pe_0_04 : BIT_VECTOR := X"178050103F4000478FFFFFFFFDEFF27740C01004C18A00067121A6803680F028";
constant pe_0_05 : BIT_VECTOR := X"A80111A8A8CEFFEF11ADF4F89A000017805D80103F4901100178050103F66000";
constant pe_0_06 : BIT_VECTOR := X"FF2FF88211C7CE922E00004A820F1FF60CFF8539776C819776A209AF6F178E01";
constant pe_0_07 : BIT_VECTOR := X"8BEFFFFFFFFF8608F08708D08F08FFC18FF7C1C7192BB7F0C1F142572F34FF8F";
constant pe_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFF1D0011FE408DEFEACE8ACE8A111048FD118BF9F";
constant pe_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_1 ----------------------------------------------------------------------------------
constant pe_1_00 : BIT_VECTOR := X"40889A8C32D8173CD0DD1FDB9742F1FEA0DA0F8003B4EDC10CBBBC3334444441";
constant pe_1_01 : BIT_VECTOR := X"45ABA3728F58889E29987F8F81811811011B07922211881886A1BEB8794F8142";
constant pe_1_02 : BIT_VECTOR := X"A24464333868037290702970F886AA04B3F4F09BB91F1D8450422391EF845042";
constant pe_1_03 : BIT_VECTOR := X"F8850B80118000E28E011A0A005A938445A5A865A86A30230A0090A821B8CA53";
constant pe_1_04 : BIT_VECTOR := X"288980E892588C880368ACE0CCD0908F4830498EEEF5836BA0058B8901780001";
constant pe_1_05 : BIT_VECTOR := X"26297A869733A86685A8061896980928898A80E892188D209288980E89238809";
constant pe_1_06 : BIT_VECTOR := X"C90233080129F0DEC120088EC29808222ECD097C240A06C68AE04444F0440D31";
constant pe_1_07 : BIT_VECTOR := X"FDDD1FDB975308908908908908908FF901D19091E0FF8233832B44242902D10D";
constant pe_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFEF986439FB0CD0CA0ECA86425AA220D934A6D00";
constant pe_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_2 ----------------------------------------------------------------------------------
constant pe_2_00 : BIT_VECTOR := X"D411EBB17F11611FF67332222222427770770F1011103F546333334444444440";
constant pe_2_01 : BIT_VECTOR := X"7F1C481F3105762E44F1AFC16864D224F04E04F0000032122040C212C0D1E0FF";
constant pe_2_02 : BIT_VECTOR := X"E4051F0EFF550E1FBC10F11016674A021AFC1001600482DF00007F1742DF0000";
constant pe_2_03 : BIT_VECTOR := X"F1240E400F8000E41D0DDC0E004EDE7AEF1F101F111E0010000000EF00050EF0";
constant pe_2_04 : BIT_VECTOR := X"08B0B0701F1080BB500000011FF6F01F12E3001DF0F13411C000D15000130004";
constant pe_2_05 : BIT_VECTOR := X"040DDDFFFF00FFF3117F012B70110008B0BF30701F101560008B0B0701F10200";
constant pe_2_06 : BIT_VECTOR := X"1F03F50B001F502AA027C1100F0361BFF1325FF75541557555F02D30F03056D4";
constant pe_2_07 : BIT_VECTOR := X"4B733222222250056050056054053F1551173616655113F533F14711FF013350";
constant pe_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFB1111F1005FF6F1104444889D31150945F124E";
constant pe_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_3 ----------------------------------------------------------------------------------
constant pe_3_00 : BIT_VECTOR := X"2F89288085C8800BBBB9999999999D0F1CF1929C999EEBE26CCCCCCCCCCCCCCC";
constant pe_3_01 : BIT_VECTOR := X"8402280580C33380F5210EF03636F3629C29CF0CCC6633633FFE2D031EF02F45";
constant pe_3_02 : BIT_VECTOR := X"2FC8D5E22499C205008C588C033F115D00EF05E00EC86D2EEC8884078D2EEC88";
constant pe_3_03 : BIT_VECTOR := X"CDEFC2FCC57CCC7F80C222C7CCF22F7124040E84088FECEEC6CC6C22FFC3F22E";
constant pe_3_04 : BIT_VECTOR := X"5EBEB0F4EEDEEEBB999999999BBBEC8CDEC21E800ECDEFD0FCCF20EECCDECECF";
constant pe_3_05 : BIT_VECTOR := X"E9D1111011DD4459FF2C9D9B2D99C45EBEBC20F4EEDEE09C45EBEB0F4EEDEEC4";
constant pe_3_06 : BIT_VECTOR := X"9EC848C2CF8F8C801C6908988FE8987FF099911F999090F999CD5537CD979F52";
constant pe_3_07 : BIT_VECTOR := X"90B9999999999EE9EE9EE9EE9EE9E40099999999F98008489858F188FEC89999";
constant pe_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFCD999940EE9BBB088888888801F89990F12099B";
constant pe_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_0 ----------------------------------------------------------------------------------
constant po_0_00 : BIT_VECTOR := X"33873F90CFE17C6CF82DFFFFFFFFF01F3DE3D8F575570D4F00FB732BDF13579B";
constant po_0_01 : BIT_VECTOR := X"7FD63A8F706911F143FFFF04121691C90A90A6A0784699C990B001011904A95F";
constant po_0_02 : BIT_VECTOR := X"AF548FEA0FF007FF7870F720791E11110FF045F00803EC1F2B617FD7FC1F2B61";
constant po_0_03 : BIT_VECTOR := X"0F060140039AE2EA01E4134A324BED8ACBFAE017C31870058A549A4018098F95";
constant po_0_04 : BIT_VECTOR := X"03F5300017805010FFFFFFFFFFF82F0610693D61D0AA06B0D0B16C0281206441";
constant po_0_05 : BIT_VECTOR := X"6F911A1919741FFE808AFFFFFC100103F1209200178059E0103F770001780501";
constant po_0_06 : BIT_VECTOR := X"FFF98FFC00199BA82FC99876971B88CABCFFF042A77AB10A7749118069306F10";
constant po_0_07 : BIT_VECTOR := X"EFADFFFFFFFFF08C08F08D08608B09D8AFFEE88D8901C40F70FD03606CF1BFFF";
constant po_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFF2232F19B9E0DF819BDF9BDF9C1127CFFC1B8FFD";
constant po_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_1 ----------------------------------------------------------------------------------
constant po_1_00 : BIT_VECTOR := X"9C88F99A23981F860F6CC0ECA863F03EB1FB0EE902A1FCD180BBBBB333444444";
constant po_1_01 : BIT_VECTOR := X"F541A4239820930F299B8688501072009EB9A1991112332653810E9286880383";
constant po_1_02 : BIT_VECTOR := X"218445A23977991398063986161EBB2094288F48BA81E5B50413F321F5B50413";
constant po_1_03 : BIT_VECTOR := X"119B1B01AA081AAE8FFA001AA3349038514749704970F2302AA1A9A8B8871852";
constant po_1_04 : BIT_VECTOR := X"8924880928898D1882479BDF1D0F689F09B0F4BFFF4B9B49888A80908AA9BAB0";
constant po_1_05 : BIT_VECTOR := X"230A8697A86BB976E22F0001E8660E8920880809288987C0E89228809288980E";
constant po_1_06 : BIT_VECTOR := X"ED89322888000EECD22190EFD138992032DECA86B350970B79BA43144CB44C33";
constant po_1_07 : BIT_VECTOR := X"D0CCC0ECA864290890890890890890EF80CC8118D8E0E1322239A5351282FC0C";
constant po_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFBE6695F2BEAE0FDB1FDB9753E402AFCE85CEECC";
constant po_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_2 ----------------------------------------------------------------------------------
constant po_2_00 : BIT_VECTOR := X"113C13B87F1F21E1E47733222222F07372172F11D1100F0E0033333444444444";
constant po_2_01 : BIT_VECTOR := X"17F0488F1100000C00DFAA114040140FD0ED0F0DD000400404220F04CE11012F";
constant po_2_02 : BIT_VECTOR := X"0E7AEF108FF55F6F1BE1F111F50048010AA11F2246FD411F0DF017F0411F0DF0";
constant po_2_03 : BIT_VECTOR := X"7F017AD7EC0DFEED3D1E00DEDCE4F0ED51F1F010F11011000EFFEDE1077046F0";
constant po_2_04 : BIT_VECTOR := X"01F1040008B0B0AFF000000011E46F510014F11DF0440140222E80007CE01ECB";
constant po_2_05 : BIT_VECTOR := X"F14DDFDFDFF00FFF4101003201000701F109430008B0B410701F1010008B0B07";
constant po_2_06 : BIT_VECTOR := X"01F77F1312605522AF34BEC10001753001322DFF555E157555073D0DF70DF139";
constant po_2_07 : BIT_VECTOR := X"F6B733222222205C05705705605504E4011136711BD4107F13F1171500FD1330";
constant po_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFB000111FF301E4D110044448F063D100951E22F";
constant po_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_3 ----------------------------------------------------------------------------------
constant po_3_00 : BIT_VECTOR := X"0C2F0E8E840F8020B99B99999999CCF309009209F99CEBEB06CCCCCCCCCCCCCC";
constant po_3_01 : BIT_VECTOR := X"085C988408CFFFC1E37C0189FCFCCFC20E20EF3EF66CFFCFFF33ECEF1089C034";
constant po_3_02 : BIT_VECTOR := X"E731240E64499F7400284088FFFC00E1E0189CDEF12F800EC2F8085C800EC2F8";
constant po_3_03 : BIT_VECTOR := X"15E01101FFF25F22310FCC222FF17C228D505E8C588C0EECE22F22F6C33FF37C";
constant po_3_04 : BIT_VECTOR := X"4EEDEEC45EBEBEBEE999999999B99E805E0FCD011E99E01EEEEF7CECEFFE0F21";
constant po_3_05 : BIT_VECTOR := X"99F11011110EE44793309999D0000F4EEDEEFBC45EBEBF30F4EEDEEC45EBEB0F";
constant po_3_06 : BIT_VECTOR := X"99E28588EE9C98880E8F02F08CC8888CC89991109992009999EF9FF52FE52091";
constant po_3_07 : BIT_VECTOR := X"BB1B999999999E9EE9EE9EE9EE9EE95F3990999902280C8588408088CCEF0999";
constant po_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFCE000905CEE0B91888888888C592F099100299B";
constant po_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

end prog_mem_content;



library IEEE;
use IEEE.STD_LOGIC_1164.all;

package prog_mem_content is

-- content of pe_0 ----------------------------------------------------------------------------------
constant pe_0_00 : BIT_VECTOR := X"E033C94222AF38FC23C40FFFFF1FF883412492595C55506EF12801ACE02468AB";
constant pe_0_01 : BIT_VECTOR := X"5077870EBC9F960558E9D4489ACC80D8D85C8E0A19F9811A081F8F068DC8002A";
constant pe_0_02 : BIT_VECTOR := X"DEF0DFFFFFFFF33C3C1B0EE8E05BC9F950CC8C805C9B0D8C91A0D6C9F9A8C9F9";
constant pe_0_03 : BIT_VECTOR := X"0071C10FEF70CF0071C1088CF071C100A90479D0F1DFE08EDF940923E5351AC1";
constant pe_0_04 : BIT_VECTOR := X"BEEA8301F08DE8AD88DD10ED8BF110FFDBEEA8501F08DE8AD8FFFF010FF592CF";
constant pe_0_05 : BIT_VECTOR := X"C269FB6CA69FB5C359FB5CB59FB4C449FB4CC49FB00CFFFF8BD10ED89F1F0FFD";
constant pe_0_06 : BIT_VECTOR := X"EE197969594939291909796959493929190080FC23B9110FF7C179FB7C979FB6";
constant pe_0_07 : BIT_VECTOR := X"9B8FFFF3C03C07C03E066E02E0C06E05C05C01C05E04E00E04E00E0CFFDAEA51";
constant pe_0_08 : BIT_VECTOR := X"0E62044FD0C210530AA0392B9B7841467CDAAE0238CDB10C8988FFFFD33422A3";
constant pe_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF08D0FF801FCEB916180B8CA5CD7129";
constant pe_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_1 ----------------------------------------------------------------------------------
constant pe_1_00 : BIT_VECTOR := X"BB1FFF333394F942AFF24C0ECA2664F3FEA0DA0F8003B4EDC100101112222221";
constant pe_1_01 : BIT_VECTOR := X"F411A366FE118F111CC6E11CEEECDCC44444555E477BE11E445A0044556AABAD";
constant pe_1_02 : BIT_VECTOR := X"CD0CCCACE0CFFF23FF2F4116344F518FF411A3EEF1D2CCFDDDFCCFD77BE6755A";
constant pe_1_03 : BIT_VECTOR := X"881EEE19C60781881EEE1889181EEE1222122E12EE0BDE2445555222422322D0";
constant pe_1_04 : BIT_VECTOR := X"18800A8F88881108D1B8088FFC88D1E8F18800E8F88881108DD1FD0EEFB81881";
constant pe_1_05 : BIT_VECTOR := X"8A98BD88A98BD88A98BD88A98BD88A98BD88A98BDB8FDF1D178088FF88881E8F";
constant pe_1_06 : BIT_VECTOR := X"CC188888888888888888888888888888888E8992AFF2888D188A98BD88A98BD8";
constant pe_1_07 : BIT_VECTOR := X"2CEFD8689AA9AA9AABB82BB2BB8AABB89AA9AA9AABB8BB8BB8BB8BBF1D16C126";
constant pe_1_08 : BIT_VECTOR := X"ED4266C5C1B95544D46252510E010733B9AFCF3F6085289B888868DF9CF8868C";
constant pe_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8083666B4B8C96E86474E1B668E9C4";
constant pe_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_2 ----------------------------------------------------------------------------------
constant pe_2_00 : BIT_VECTOR := X"F07F1F77751D43F1FF1F033222D2C5417770770F1011102F54CC204444444440";
constant pe_2_01 : BIT_VECTOR := X"1176E63510FF11176EE1576F11E11FDFF3711F010FF11761F191FF371F1FFF51";
constant pe_2_02 : BIT_VECTOR := X"FF6C7300011E5471F1F1176F63711F111176E63F11F63711EC03711FF1111FF1";
constant pe_2_03 : BIT_VECTOR := X"11DFFB0F14203F11DFFA0303F1DFF00D99CBB721472F11B77667777664766516";
constant pe_2_04 : BIT_VECTOR := X"7557F1F657755F5D471D7752E1D7170503553F1F657355F1D0332207003B433F";
constant pe_2_05 : BIT_VECTOR := X"1957F131917F171957F131917F171957F131917F1111001171D7756E1D717454";
constant pe_2_06 : BIT_VECTOR := X"11075757575757575757171717171717171630F1FF1F0113371957F131917F17";
constant pe_2_07 : BIT_VECTOR := X"01E222231F11F11F5F073F03F01F1F071F51F51F1F07F07F03F03F0111F010FF";
constant pe_2_08 : BIT_VECTOR := X"2EEA1D77CF6D3C9DFCBC13BE3726785FD449271BC59B2001F7F3000091F1AAE1";
constant pe_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB0102C549615E98153EDD68A658536";
constant pe_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_3 ----------------------------------------------------------------------------------
constant pe_3_00 : BIT_VECTOR := X"4E91019229029F590102E9999907269D0F1CF1929C999EEBE22501CCCCCCCCCC";
constant pe_3_01 : BIT_VECTOR := X"08990982091400899000299000298520582984E0514009905800058284907790";
constant pe_3_02 : BIT_VECTOR := X"BBB5B999999C19291050899098209100089909820919820911E8209140089140";
constant pe_3_03 : BIT_VECTOR := X"88F00EE405DEF588F00EEE3F58F00EEBBBBBBF9E5F940E888EEEEEEEEEEEE909";
constant pe_3_04 : BIT_VECTOR := X"82282D222282228282D222282D22D282882282D2222822282899990F4EEBFBF5";
constant pe_3_05 : BIT_VECTOR := X"958240895824089582408958240895824089582400E099992D222282D22D2828";
constant pe_3_06 : BIT_VECTOR := X"00E28282828282828282828282828282828EFE590102E1999895824089582408";
constant pe_3_07 : BIT_VECTOR := X"D02999989589589584E884E84E9584E89589589584E84E84E84E84E099DE03D2";
constant pe_3_08 : BIT_VECTOR := X"35E285A90FB9A3F4E4CFDE368219CDA3FAD58D0679B90EE00202999900C90120";
constant pe_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF110372659EA51DFC303BDA775DC9D0";
constant pe_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_0 ----------------------------------------------------------------------------------
constant po_0_00 : BIT_VECTOR := X"C0CF20890020DF003B20BFFFFFAC0CF0173DE3D8F575570D4F02B00BDF13579B";
constant po_0_01 : BIT_VECTOR := X"06AC9F980668A0E8C91580C948D33E09F9B22A081F8E85C8E0A29F957A09AA21";
constant po_0_02 : BIT_VECTOR := X"EF81EF8FFFFF8A08F2F056C9F980DD8D01AC9F910BB8960AA8F9B09987878888";
constant po_0_03 : BIT_VECTOR := X"87A1D0DCFFE08047A1D0D2920AA1D0BEE8310FAFFEA1F20FBCBA98FEDCBA99D0";
constant po_0_04 : BIT_VECTOR := X"C8CD10E98AF100BF9FEEE8401F0CDE8EDC8ED10E98CF120BF9CFFFD0012804C0";
constant po_0_05 : BIT_VECTOR := X"9FB2C629FB2CE29FB1C719FB1CF19FB0C809FB0C01808FFFFEEE8201F0CDE8ED";
constant po_0_06 : BIT_VECTOR := X"428FFEEDDCCBBAA9988FFEEDDCCBBAA99880B0103A204EBCF89FB3C539FB3CD3";
constant po_0_07 : BIT_VECTOR := X"838BFFF87E03E07E0C072C06C02E0C021E05E01E0C01C04C00C04C008F0E80FE";
constant po_0_08 : BIT_VECTOR := X"AB80F9E433A80F23A8E10F6AC205315732279B7F721E808088B48FFF1C81C2FC";
constant po_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6020C0CBD2987E8D765B445E4E74C4";
constant po_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_1 ----------------------------------------------------------------------------------
constant po_1_00 : BIT_VECTOR := X"7AADEDEF2325FF42BDE30D1FDB0626F03EB1FB0EE902A1FCD180280111222222";
constant po_1_01 : BIT_VECTOR := X"44F6B5FF6110011FEDDEEEDD2EE11DD55AE11E445A66444555E411844E4BBBB1";
constant po_1_02 : BIT_VECTOR := X"C0FDDD0BDF1D0F221E344F57BFF4110344F1B5FE011CEFC11CC6FC1166661144";
constant po_1_03 : BIT_VECTOR := X"28FFFF0287B86148FFFF057815FFFF052221222DFF20AF234555522242232E12";
constant po_1_04 : BIT_VECTOR := X"D198088FFA88B1E8F18800C8F88881108D1D8088FFE88F1E8FEC0EB0FBE98891";
constant po_1_05 : BIT_VECTOR := X"8BD88A98BD88A98BD88A98BD88A98BD88A98BD88A1690E0C1880088F88881108";
constant po_1_06 : BIT_VECTOR := X"91089898989898989898989898989898989FE902BDE3602AC08BD88A98BD88A9";
constant po_1_07 : BIT_VECTOR := X"A0A6EC709BB9BB9BB8AA92AA2AABB9AA9BB9BB9BB8AA8AA8AA8AA8AA0C8C0B1C";
constant po_1_08 : BIT_VECTOR := X"30B941741FD34903A5BB02D52B8023EF97A4CA667D8F0828009207CE08A8F723";
constant po_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3203626B248288915FB87B2AF43EA2";
constant po_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_2 ----------------------------------------------------------------------------------
constant po_2_00 : BIT_VECTOR := X"1F11F0F1FF500413F1F0033222047CF07372172F11D1100F0E0B010444444444";
constant po_2_01 : BIT_VECTOR := X"3711E111176FF3510EC0310F62676F0FF11761F191FF3711F010FF17F1EF7757";
constant po_2_02 : BIT_VECTOR := X"1E497350001100316FF3711F111176F63711E117176F11176EE11176FF3776FF";
constant po_2_03 : BIT_VECTOR := X"2B5DF0015F10812B5DF00253225DF002013AFF51F1505017477777333333372A";
constant po_2_04 : BIT_VECTOR := X"471D7756E1D7174543553F1F657355F1D071D7752E1D7170501332F0004BF011";
constant po_2_05 : BIT_VECTOR := X"7F171957F131917F171957F131917F171957F131A4F150117557F1F657755F5D";
constant po_2_06 : BIT_VECTOR := X"E007575757575757575313131313131313101103F1F00021357F171957F13191";
constant po_2_07 : BIT_VECTOR := X"D0F122253F07F07F01F571F51F5F01F17F03F03F01F11F51F51F11F1510103F1";
constant po_2_08 : BIT_VECTOR := X"AB48C3D7C215F8F5BF9BD430A52A351C60F0D6B5BB0F53C65514500079D11AF1";
constant po_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF04047C6F8DF941E9E6AF6E8A9D92C";
constant po_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_3 ----------------------------------------------------------------------------------
constant po_3_00 : BIT_VECTOR := X"95900800779EC238100EC999990656CCF309009209F99CEBEB02006CCCCCCCCC";
constant po_3_01 : BIT_VECTOR := X"8209100089905820911E8891982994E140099058000582984E05140220512299";
constant po_3_02 : BIT_VECTOR := X"0B90B9999999FE88904820910008990982091002899000899000089905829905";
constant po_3_03 : BIT_VECTOR := X"DB911ECD540EE3DB911ECDFB3D911ECDEEEBEE9040995EE8E888888888888F9E";
constant po_3_04 : BIT_VECTOR := X"82D222282D22D282882282D222282228282D222282D22D28280999CC45EBE3B3";
constant po_3_05 : BIT_VECTOR := X"24089582408958240895824089582408958240895298999982282D2222822282";
constant po_3_06 : BIT_VECTOR := X"DDC88888888888888888888888888888888E03C8100ECC009924089582408958";
constant po_3_07 : BIT_VECTOR := X"2C20999984E84E84E95889589584E95884E84E84E95895895895895899E0DF50";
constant po_3_08 : BIT_VECTOR := X"0D18D731ED2F8A78FC35E8BA17E9C1FC2CAF772C7CEC99DE99EF9999912100E0";
constant po_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4036761060DE919B0681C20EA6765";
constant po_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

end prog_mem_content;



library IEEE;
use IEEE.STD_LOGIC_1164.all;

package prog_mem_content is

-- content of pe_0 ----------------------------------------------------------------------------------
constant pe_0_00 : BIT_VECTOR := X"873F90CFE17C6CF82DFFFFFFFF048B412492595C5550AEF10B73F9468ACE024F";
constant pe_0_01 : BIT_VECTOR := X"D63A8F706911F143FFFF04121691C90A90A6A0784699C990B001011904A95F33";
constant pe_0_02 : BIT_VECTOR := X"548FEA0FF007FF7870F720791E11110FF045600803EC1F2B617FD7FC1F2B617F";
constant pe_0_03 : BIT_VECTOR := X"060140039AE2EA01E4134A324BED8AC1FAE017C31870058A549A4018098F95AF";
constant pe_0_04 : BIT_VECTOR := X"A1919741FFE808AFFFFFFFFFF82F0610693461D0AA06B0D0B16C02812064410F";
constant pe_0_05 : BIT_VECTOR := X"A7050017805F0103FC3050017805F50F042A77AB10A7749118069306F106F911";
constant pe_0_06 : BIT_VECTOR := X"608F08708D08F08FFC18FF7C1C7192BB7F0C1F142572F34FF7F0104FFF00103F";
constant pe_0_07 : BIT_VECTOR := X"FFFFFFFFFFFF160011FE308DEFEACE8ACE8A111048FD118BF9F8BEFFFFFFFFF8";
constant pe_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_1 ----------------------------------------------------------------------------------
constant pe_1_00 : BIT_VECTOR := X"88F99A23981F860F6CC0ECA86307F7FEA0DA0F8003B4EDC1055546DDDDDDEEE1";
constant pe_1_01 : BIT_VECTOR := X"41A4239820930F299B8688501072009EB9A1991112332653810E92868803839C";
constant pe_1_02 : BIT_VECTOR := X"8445A23977991398063986161EBB2094288FE8BA81E5B50413F321F5B50413F5";
constant pe_1_03 : BIT_VECTOR := X"9B1B01AA081AAE8FFA001AA33490385A4749704970F2302AA1A9A8B887185221";
constant pe_1_04 : BIT_VECTOR := X"697A86BB976E22F2479BDF1D0F689F09B0FEBFFF4B9B49888A80908AA9BAB011";
constant pe_1_05 : BIT_VECTOR := X"5888092889880E892788809288988888A86B350970B79BA43144CB44C33230A8";
constant pe_1_06 : BIT_VECTOR := X"8908908908908908FF901D19091E0FF8233832B44242902D1A00E8928A90E892";
constant pe_1_07 : BIT_VECTOR := X"FFFFFFFFFFFFE6986439FB0CD0CA0ECA86425AA220D934A6D00FDDD1FDB97530";
constant pe_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_2 ----------------------------------------------------------------------------------
constant pe_2_00 : BIT_VECTOR := X"3C13B87F1F21E1E47733222222F5427770770F1011103F546333333333333330";
constant pe_2_01 : BIT_VECTOR := X"F0488F1100000C00DFAA114040140FD0ED0F0DD000400404220F04CE11012F11";
constant pe_2_02 : BIT_VECTOR := X"7AEF108FF55F6F1BE1F111F50048010AA11F1246FD411F0DF017F0411F0DF017";
constant pe_2_03 : BIT_VECTOR := X"017AD7EC0DFEED3D1E00DEDCE4F0ED50F1F010F11011000EFFEDE1077046F00E";
constant pe_2_04 : BIT_VECTOR := X"FDFDFF00FFF4101000000011E46F510014F01DF0440140222E80007CE01ECB7F";
constant pe_2_05 : BIT_VECTOR := X"00130008B0B00701F00430008B0B03FFDFF555E157555073D0DF70DF139F14DD";
constant pe_2_06 : BIT_VECTOR := X"0056050056054053F1551173616655113F533F14711FF0133F00700F3300701F";
constant pe_2_07 : BIT_VECTOR := X"FFFFFFFFFFFFFC1111F1005FF6F1104444889D31150945F124E4B73322222225";
constant pe_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_3 ----------------------------------------------------------------------------------
constant pe_3_00 : BIT_VECTOR := X"2F0E8E840F8020B99B99999999F69D0F1CF1929C999EEBE26CCCCCCCCCCCCCCC";
constant pe_3_01 : BIT_VECTOR := X"5C988408CFFFC1E37C0189FCFCCFC20E20EF3EF66CFFCFFF33ECEF1089C0340C";
constant pe_3_02 : BIT_VECTOR := X"31240E64499F7400284088FFFC00E1E0189CDEF12F800EC2F8085C800EC2F808";
constant pe_3_03 : BIT_VECTOR := X"E01101FFF25F22310FCC222FF17C228D505E8C588C0EECE22F22F6C33FF37CE7";
constant pe_3_04 : BIT_VECTOR := X"011110EE4479330999999999B99E805E0FCD011E99E01EEEEF7CECEFFE0F2115";
constant pe_3_05 : BIT_VECTOR := X"DE6BC45EBEB70F4EEDE6BC45EBEB7BEE1109992009999EF9FF52FE5209199F11";
constant pe_3_06 : BIT_VECTOR := X"EE9EE9EE9EE9EE9E40099999999F98008489858F188FEC899C90F4EE99E0F4EE";
constant pe_3_07 : BIT_VECTOR := X"FFFFFFFFFFFFCD999940EE9BBB088888888801F89990F12099B90B9999999999";
constant pe_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_0 ----------------------------------------------------------------------------------
constant po_0_00 : BIT_VECTOR := X"9049A89DFA409ADEFEFFFFFFFFF3F01F3DE3D8F575570D4F00951DC579BDF135";
constant po_0_01 : BIT_VECTOR := X"F71A99E97F333928581FF7380C06E01E31A688913210D0309001565127949FF8";
constant po_0_02 : BIT_VECTOR := X"99C8F031F10A19E9019C318794912196FF7110690BF054F0320EF7FED4F0320E";
constant po_0_03 : BIT_VECTOR := X"D08D0060F64589104EB435E9B8936F58FEF700F7207220066A94D85196815101";
constant po_0_04 : BIT_VECTOR := X"11A8A8CEFFEF11A8FFFFFFFFDEFF277B0C01004C18100767121A68036F0F0288";
constant po_0_05 : BIT_VECTOR := X"805F0103FB6050017805F0103FD005478539776C819776A209AF6F178E01A801";
constant po_0_06 : BIT_VECTOR := X"08C08F08D08608B09D8AFFEE88D8901C40F70FD03606CF1BFFFF00113F000017";
constant po_0_07 : BIT_VECTOR := X"FFFFFFFFFFFF8232F19B980DF819BDF9BDF9C1127CFFC1B8FFDEFADFFFFFFFFF";
constant po_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_1 ----------------------------------------------------------------------------------
constant po_1_00 : BIT_VECTOR := X"0889A8C32D8173CD0DD1FDB97427F03EB1FB0EE902A1FCD18055544DDDDDDEEE";
constant po_1_01 : BIT_VECTOR := X"5ABA3728F58889E29987F8F81811811011B07922211881886A1B8B8794F81424";
constant po_1_02 : BIT_VECTOR := X"244E4333868037290702970F886AA0DB3F4F09BB91F178450422391E88450424";
constant po_1_03 : BIT_VECTOR := X"1850B80118000E28E011A0A005A938445A5A865A86A30230A0090A821B8CA53A";
constant po_1_04 : BIT_VECTOR := X"7A869733A86685A0368ACE0CCD0908FD830498EEEFF83FBA0058B8901080001F";
constant po_1_05 : BIT_VECTOR := X"89880E8926888092889880E892888888097C240A06C68AE04444F0440D312629";
constant po_1_06 : BIT_VECTOR := X"90890890890890890EF80CC8118D8E0E1322239A5351282FC0000928C9A80928";
constant po_1_07 : BIT_VECTOR := X"FFFFFFFFFFFF1E6695F2BEAE0FDB1FDB9753E402AFCE85CEECCD0CCC0ECA8642";
constant po_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_2 ----------------------------------------------------------------------------------
constant po_2_00 : BIT_VECTOR := X"411EBB17F11611FF673322222224F07372172F11D1100F0E0033333333333333";
constant po_2_01 : BIT_VECTOR := X"F1C481F3105762E44F1AFC16864D224F04E04F0000032122040C212C0D1E0FFD";
constant po_2_02 : BIT_VECTOR := X"4050F0EFF550E1FBC10F11016674A011AFC1001600482DF00007F1742DF00007";
constant po_2_03 : BIT_VECTOR := X"1240E400F8000E41D0DDC0E004EDE7AEF1F101F111E0010000000EF00050EF0E";
constant po_2_04 : BIT_VECTOR := X"DDFFFF00FFF3117500000011FF6F01F02E3001DF0F03401C000D15000130004F";
constant po_2_05 : BIT_VECTOR := X"B0B00701F00230008B0B00701F0083BB5FF75541557555F02D30F03056D4040D";
constant po_2_06 : BIT_VECTOR := X"05C05705705605504E4011136711BD4107F13F1171500FD13300000E03090008";
constant po_2_07 : BIT_VECTOR := X"FFFFFFFFFFFFC000111FFD01E4D110044448F063D100951E22FF6B7332222222";
constant po_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_3 ----------------------------------------------------------------------------------
constant po_3_00 : BIT_VECTOR := X"F89288085C8800BBBB9999999997CCF309009209F99CEBEB06CCCCCCCCCCCCCC";
constant po_3_01 : BIT_VECTOR := X"402280580C33380F5210EF03636F3629C29CF0CCC6633633FFE2D031EF02F452";
constant po_3_02 : BIT_VECTOR := X"FC8D5E22499C205008C588C033F115D00EF05E00EC86D2EEC8884078D2EEC888";
constant po_3_03 : BIT_VECTOR := X"DEFC2FCC57CCC7F80C222C7CCF22F7124040E84088FECEEC6CC6C22FFC3F22E2";
constant po_3_04 : BIT_VECTOR := X"111011DD4459FF2999999999BBBEC8CDEC21E800ECDEFD0FCCF20EECCDECECFC";
constant po_3_05 : BIT_VECTOR := X"BEB70F4EEDE6BC45EBEB70F4EEDE6BBB911F999090F999CD5537CD979F52E9D1";
constant po_3_06 : BIT_VECTOR := X"E9EE9EE9EE9EE9EE95F3990999902280C8588408088CCEF09999C45ED9EEC45E";
constant po_3_07 : BIT_VECTOR := X"FFFFFFFFFFFFCE000905CEE0B91888888888C592F099100299BBB1B999999999";
constant po_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

end prog_mem_content;


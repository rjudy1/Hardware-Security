
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package prog_mem_content is

-- content of pe_0 ----------------------------------------------------------------------------------
constant pe_0_00 : BIT_VECTOR := X"95F33873F90CFE17C6CF82DFFFFFFFF048B412492595C55506EF1002468ACE05";
constant pe_0_01 : BIT_VECTOR := X"B617FD63A8F706911F143FFFF04121691C90A90A6A0784699C990B001011904A";
constant pe_0_02 : BIT_VECTOR := X"F95AF548FEA0FF007FF7870F720791E11110FF045400803EC1F2B617FD7FC1F2";
constant pe_0_03 : BIT_VECTOR := X"4410F060140039AE2EA01E4134A324BED8AC1FAE017C31870058A549A4018098";
constant pe_0_04 : BIT_VECTOR := X"6F911A1919741FFE808AFFFFFFFFFF82F0610693261D0AA06B0D0B16C0281206";
constant pe_0_05 : BIT_VECTOR := X"F0C001485F010EF205001485F010EF805950F042A77AB10A7749118069306F10";
constant pe_0_06 : BIT_VECTOR := X"1048FD118BF9F8BEFFFFFFFFF8FF7C1C7192BB7F0C1F142572F34FF9001182FE";
constant pe_0_07 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF100011FE308DEFEACE8ACE8A11";
constant pe_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_1 ----------------------------------------------------------------------------------
constant pe_1_00 : BIT_VECTOR := X"3839C88F99A23981F860F6CC0ECA86307F7FEA0DA0F8003B4EDC10AAAAAAAAB1";
constant pe_1_01 : BIT_VECTOR := X"413F541A4239820930F299B8688501072009EB9A1991112332653810E9286880";
constant pe_1_02 : BIT_VECTOR := X"852218445A23977991398063986161EBB2094288FE8BA81E5B50413F321F5B50";
constant pe_1_03 : BIT_VECTOR := X"AB0119B1B01AA081AAE8FFA001AA33490385A4749704970F2302AA1A9A8B8871";
constant pe_1_04 : BIT_VECTOR := X"230A8697A86BB976E22F2479BDF1D0F689F09B0FEBFFF4B9B49888A80908AA9B";
constant pe_1_05 : BIT_VECTOR := X"9A809288880E89288809288880E8928880888A86B350970B79BA43144CB44C33";
constant pe_1_06 : BIT_VECTOR := X"A220D934A6D00FDDD1FDB975301D19091E0FF8233832B44242902D1A09288009";
constant pe_1_07 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE9986439FB0CD0CA0ECA86425A";
constant pe_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_2 ----------------------------------------------------------------------------------
constant pe_2_00 : BIT_VECTOR := X"12F113C13B87F1F21E1E47733222222F5427770770F1011102F5463333333330";
constant pe_2_01 : BIT_VECTOR := X"DF017F0488F1100000C00DFAA114040140FD0ED0F0DD000400404220F04CE110";
constant pe_2_02 : BIT_VECTOR := X"6F00E7AEF108FF55F6F1BE1F111F50048010AA11F1246FD411F0DF017F0411F0";
constant pe_2_03 : BIT_VECTOR := X"ECB7F017AD7EC0DFEED3D1E00DEDCE4F0ED50F1F010F11011000EFFEDE107704";
constant pe_2_04 : BIT_VECTOR := X"F14DDFDFDFF00FFF4101000000011E46F510014F01DF0440140222E80007CE01";
constant pe_2_05 : BIT_VECTOR := X"3070008BB0070172230008BB00701788343FFDFF555E157555073D0DF70DF139";
constant pe_2_06 : BIT_VECTOR := X"31150945F124E4B733222222251173616655113F533F14711FF0133F000AB000";
constant pe_2_07 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1111F1005FF6F1104444889D";
constant pe_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_3 ----------------------------------------------------------------------------------
constant pe_3_00 : BIT_VECTOR := X"0340C2F0E8E840F8020B99B99999999F69D0F1CF1929C999EEBE26CCCCCCCCCC";
constant pe_3_01 : BIT_VECTOR := X"2F8085C988408CFFFC1E37C0189FCFCCFC20E20EF3EF66CFFCFFF33ECEF1089C";
constant pe_3_02 : BIT_VECTOR := X"37CE731240E64499F7400284088FFFC00E1E0189CDEF12F800EC2F8085C800EC";
constant pe_3_03 : BIT_VECTOR := X"F2115E01101FFF25F22310FCC222FF17C228D505E8C588C0EECE22F22F6C33FF";
constant pe_3_04 : BIT_VECTOR := X"99F11011110EE4479330999999999B99E805E0FCD011E99E01EEEEF7CECEFFE0";
constant pe_3_05 : BIT_VECTOR := X"9EEC45EBB70F4EEE6BC45EBB70F4EEE6BFBEE1109992009999EF9FF52FE52091";
constant pe_3_06 : BIT_VECTOR := X"F89990F12099B90B99999999999999999F98008489858F188FEC899CC45EBC9D";
constant pe_3_07 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCD999940EE9BBB088888888801";
constant pe_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_0 ----------------------------------------------------------------------------------
constant po_0_00 : BIT_VECTOR := X"49FF89049A89DFA409ADEFEFFFFFFFFF3F01B3DE3D8F575570D4F0013579BDF1";
constant po_0_01 : BIT_VECTOR := X"0320EF71A99E97F333928581FF7380C06E01E31A688913210D03090013651279";
constant po_0_02 : BIT_VECTOR := X"1510199C8F031F10A19E9019C318794912176FF7110690BF0B4F0320EF7FE34F";
constant po_0_03 : BIT_VECTOR := X"F0288B08D0060F64589104EB435E9B8936F58FEF700F7207220066A94D851968";
constant po_0_04 : BIT_VECTOR := X"1A80111A8A8CEFFEF11A8FFFFFFFFDEFF27790C01004C18F00567121A68036D0";
constant po_0_05 : BIT_VECTOR := X"FF0010EF105001485F010EF405001485F78478539776C819776A209AF6F178E0";
constant po_0_06 : BIT_VECTOR := X"127CFFC1B8FFDEFADFFFFFFFFFFFEE88D8901C40F70FD03606CF1BFF0107FFFF";
constant po_0_07 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC232F19B940DF819BDF9BDF9C1";
constant po_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_1 ----------------------------------------------------------------------------------
constant po_1_00 : BIT_VECTOR := X"814240889A8C32D8173CD0DD1FDB97427F03EB1FB0EE902A1FCD180AAAAAAAAB";
constant po_1_01 : BIT_VECTOR := X"504245ABA3728F58889E29987F8F81811811011B07922211881886A1B8B8794F";
constant po_1_02 : BIT_VECTOR := X"CA53A244E4333868037290702970F886AA0DB3F4F09BB91F148450422391E684";
constant po_1_03 : BIT_VECTOR := X"0001F1850B80118000E28E011A0A005A938445A5A865A86A30230A0090A821B8";
constant po_1_04 : BIT_VECTOR := X"126297A869733A86685A0368ACE0CCD0908FD830498EEEFE83FBA0058B890108";
constant po_1_05 : BIT_VECTOR := X"8A90E89288809288880E89288809288884888097C240A06C68AE04444F0440D3";
constant po_1_06 : BIT_VECTOR := X"02AFCE85CEECCD0CCC0ECA86420CC8118D8E0E1322239A5351282FC00E892800";
constant po_1_07 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4E6695F2BEAE0FDB1FDB9753E4";
constant po_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_2 ----------------------------------------------------------------------------------
constant po_2_00 : BIT_VECTOR := X"E0FFD411EBB17F11611FF673322222224F07272172F11D1100F0E00333333333";
constant po_2_01 : BIT_VECTOR := X"00007F1C481F3105762E44F1AFC16864D224F04E04F0000032122040C212C0D1";
constant po_2_02 : BIT_VECTOR := X"0EF0E4050F0EFF550E1FBC10F11016674A011AFC1001600482DF00007F1742DF";
constant po_2_03 : BIT_VECTOR := X"0004F1240E400F8000E41D0DDC0E004EDE7AEF1F101F111E0010000000EF0005";
constant po_2_04 : BIT_VECTOR := X"4040DDDFFFF00FFF3117500000011FF6F01F02E3001DF0F03401C000D1500013";
constant po_2_05 : BIT_VECTOR := X"330070171130008BB0070174430008BB003BB5FF75541557555F02D30F03056D";
constant po_2_06 : BIT_VECTOR := X"63D100951E22FF6B733222222211136711BD4107F13F1171500FD13307001700";
constant po_2_07 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000111FFA01E4D110044448F0";
constant po_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_3 ----------------------------------------------------------------------------------
constant po_3_00 : BIT_VECTOR := X"2F452F89288085C8800BBBB9999999997CCF309009209F99CEBEB06CCCCCCCCC";
constant po_3_01 : BIT_VECTOR := X"EC888402280580C33380F5210EF03636F3629C29CF0CCC6633633FFE2D031EF0";
constant po_3_02 : BIT_VECTOR := X"F22E2FC8D5E22499C205008C588C033F115D00EF05E00EC86D2EEC8884078D2E";
constant po_3_03 : BIT_VECTOR := X"CECFCDEFC2FCC57CCC7F80C222C7CCF22F7124040E84088FECEEC6CC6C22FFC3";
constant po_3_04 : BIT_VECTOR := X"2E9D1111011DD4459FF2999999999BBBEC8CDEC21E800ECDEFD0FCCF20EECCDE";
constant po_3_05 : BIT_VECTOR := X"99E0F4EEE6BC45EBB70F4EEE6BC45EBB7C2BB911F999090F999CD5537CD979F5";
constant po_3_06 : BIT_VECTOR := X"92F099100299BBB1B999999999990999902280C8588408088CCEF0990F4EEE99";
constant po_3_07 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCE000905CEE0B91888888888C5";
constant po_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

end prog_mem_content;



library IEEE;
use IEEE.STD_LOGIC_1164.all;

package prog_mem_content is

-- content of pe_0 ----------------------------------------------------------------------------------
constant pe_0_00 : BIT_VECTOR := X"9049A89DFA409ADEFEFFFFFFFFF88C412492595C5550AEF102EA60BDF13579BF";
constant pe_0_01 : BIT_VECTOR := X"F71A99E97F333928581FF7380C06E01E31A688913210D0309001D65127949FF8";
constant pe_0_02 : BIT_VECTOR := X"99CDF031F10A19E9019C318794912116FF7110690BF0D4F0320EF7FE54F0320E";
constant pe_0_03 : BIT_VECTOR := X"508D0060F64589104EB435E9B8936F58FEF700F7207220066A94D85196815101";
constant pe_0_04 : BIT_VECTOR := X"178050103F500478FFFFFFFFDEFF27730C01004C18900F67121A6803670F0288";
constant pe_0_05 : BIT_VECTOR := X"069306F106F911A1919741FFE808AFFFF0920000178059200178050103F76000";
constant pe_0_06 : BIT_VECTOR := X"8F08D08608B09D8AFFEE88D8901C40F70FD03606CF1BFF042A77AB10A7749118";
constant pe_0_07 : BIT_VECTOR := X"FFFFFFFF1232F19B9F0DF819BDF9BDF9C1127CFFC1B8FFDEFADFFFFFFFFF08C0";
constant pe_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_1 ----------------------------------------------------------------------------------
constant pe_1_00 : BIT_VECTOR := X"0889A8C32D8173CD0DD1FDB97426F1FEA0DA0F8003B4EDC1065557DDDEEEEEE1";
constant pe_1_01 : BIT_VECTOR := X"5ABA3728F58889E29987F8F81811811011B07922211881886A1B8B8794F81424";
constant pe_1_02 : BIT_VECTOR := X"24444333868037290702970F886AA0EB3F4F09BB91F178450422391E98450424";
constant pe_1_03 : BIT_VECTOR := X"2850B80118000E28E011A0A005A938445A5A865A86A30230A0090A821B8CA53A";
constant pe_1_04 : BIT_VECTOR := X"288980E892F88880368ACE0CCD0908FE830498EEEFF83FBA0058B8901180001F";
constant pe_1_05 : BIT_VECTOR := X"44CB44C33230A8697A86BB976E22F008A9687609288980809288980E892D8809";
constant pe_1_06 : BIT_VECTOR := X"0890890890890EF80CC8118D8E0E1322239A5351282FC0A86B350970B79BA431";
constant pe_1_07 : BIT_VECTOR := X"FFFFFFFF1E6695F2BEAE0FDB1FDB9753E402AFCE85CEECCD0CCC0ECA86429089";
constant pe_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_2 ----------------------------------------------------------------------------------
constant pe_2_00 : BIT_VECTOR := X"411EBB17F11611FF673322222229427770770F1011103F546333333333333330";
constant pe_2_01 : BIT_VECTOR := X"F1C481F3105762E44F1AFC16864D224F04E04F0000032122040C212C0D1E0FFD";
constant pe_2_02 : BIT_VECTOR := X"4051F0EFF550E1FBC10F11016674A011AFC1001600482DF00007F1742DF00007";
constant pe_2_03 : BIT_VECTOR := X"1240E400F8000E41D0DDC0E004EDE7AEF1F101F111E0010000000EF00050EF0E";
constant pe_2_04 : BIT_VECTOR := X"08B0B0701F008BB500000011FF6F01F02E3001DF0F03401C000D15000130004F";
constant pe_2_05 : BIT_VECTOR := X"DF70DF139F14DDFDFDFF00FFF41010033006110008B0B230008B0B0701F00200";
constant pe_2_06 : BIT_VECTOR := X"5705705605504E4011136711BD4107F13F1171500FD133DFF555E157555073D0";
constant pe_2_07 : BIT_VECTOR := X"FFFFFFFFC000111FFD01E4D110044448F063D100951E22FF6B733222222205C0";
constant pe_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_3 ----------------------------------------------------------------------------------
constant pe_3_00 : BIT_VECTOR := X"F89288085C8800BBBB99999999969D0F1CF1929C999EEBE26CCCCCCCCCCCCCCC";
constant pe_3_01 : BIT_VECTOR := X"402280580C33380F5210EF03636F3629C29CF0CCC6633633FFE2D031EF02F452";
constant pe_3_02 : BIT_VECTOR := X"FC8D5E22499C205008C588C033F115D00EF05E00EC86D2EEC8884078D2EEC888";
constant pe_3_03 : BIT_VECTOR := X"DEFC2FCC57CCC7F80C222C7CCF22F7124040E84088FECEEC6CC6C22FFC3F22E2";
constant pe_3_04 : BIT_VECTOR := X"5EBEB0F4EEDEEBB999999999BBBEC8CDEC21E800ECDEFD0FCCF20EECCDECECFC";
constant pe_3_05 : BIT_VECTOR := X"52FE5209199F11011110EE44793309999EDE99C45EBEBFBC45EBEB0F4EEDEEC4";
constant pe_3_06 : BIT_VECTOR := X"9EE9EE9EE9EE95F3990999902280C8588408088CCEF0991109992009999EF9FF";
constant pe_3_07 : BIT_VECTOR := X"FFFFFFFFCE000905CEE0B91888888888C592F099100299BBB1B999999999E9EE";
constant pe_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_0 ----------------------------------------------------------------------------------
constant po_0_00 : BIT_VECTOR := X"3873F90CFE17C6CF82DFFFFFFFF0F01F3DE3D8F575570D4F000C843CE02468AC";
constant po_0_01 : BIT_VECTOR := X"FD63A8F706911F143FFFF04121691C90A90A6A0784699C990B001011904A95F3";
constant po_0_02 : BIT_VECTOR := X"F548FEA0FF007FF7870F720791E11110FF045E00803EC1F2B617FD7FC1F2B617";
constant po_0_03 : BIT_VECTOR := X"F060140039AE2EA01E4134A324BED8AC6FAE017C31870058A549A4018098F95A";
constant po_0_04 : BIT_VECTOR := X"03F630001780510FFFFFFFFFFF82F0610693C61D0AA06B0D0B16C02812064410";
constant po_0_05 : BIT_VECTOR := X"AF6F178E01A80111A8A8CEFFEF11A0F8F000320103F62080103F870001780501";
constant po_0_06 : BIT_VECTOR := X"F08708D08F08FFC18FF7C1C7192BB7F0C1F142572F34FF8539776C819776A209";
constant po_0_07 : BIT_VECTOR := X"FFFFFFFFF1E0011FE308DEFEACE8ACE8A111048FD118BF9F8BEFFFFFFFFF8608";
constant po_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_1 ----------------------------------------------------------------------------------
constant po_1_00 : BIT_VECTOR := X"C88F99A23981F860F6CC0ECA8630F03EB1FB0EE902A1FCD18065555DDEEEEEEE";
constant po_1_01 : BIT_VECTOR := X"541A4239820930F299B8688501072009EB9A1991112332653810E92868803839";
constant po_1_02 : BIT_VECTOR := X"18445A23977991398063986161EBB2094288FE8BA81E5B50413F321F5B50413F";
constant po_1_03 : BIT_VECTOR := X"19B1B01AA081AAE8FFA001AA3349038504749704970F2302AA1A9A8B88718522";
constant po_1_04 : BIT_VECTOR := X"892E8809288981882479BDF1D0F689F09B0FEBFFF4B9B49888A80908AA9BAB01";
constant po_1_05 : BIT_VECTOR := X"44F0440D3126297A869733A86685AA019A89660E892B8880E892C8809288980E";
constant po_1_06 : BIT_VECTOR := X"8908908908908FF901D19091E0FF8233832B44242902D1097C240A06C68AE044";
constant po_1_07 : BIT_VECTOR := X"FFFFFFFFFE5986439FB0CD0CA0ECA86425AA220D934A6D00FDDD1FDB97530890";
constant po_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_2 ----------------------------------------------------------------------------------
constant po_2_00 : BIT_VECTOR := X"13C13B87F1F21E1E47733222222FF07372172F11D1100F0E0033333333333333";
constant po_2_01 : BIT_VECTOR := X"7F0488F1100000C00DFAA114040140FD0ED0F0DD000400404220F04CE11012F1";
constant po_2_02 : BIT_VECTOR := X"E7AEF108FF55F6F1BE1F111F50048010AA11F1246FD411F0DF017F0411F0DF01";
constant po_2_03 : BIT_VECTOR := X"F017AD7EC0DFEED3D1E00DEDCE4F0ED51F1F010F11011000EFFEDE1077046F00";
constant po_2_04 : BIT_VECTOR := X"01F0040008B0BAFF000000011E46F510014F01DF0440140222E80007CE01ECB7";
constant po_2_05 : BIT_VECTOR := X"30F03056D4040DDDFFFF00FFF3117F013090000701F00930701F0010008B0B07";
constant po_2_06 : BIT_VECTOR := X"6050056054053F1551173616655113F533F14711FF01335FF75541557555F02D";
constant po_2_07 : BIT_VECTOR := X"FFFFFFFFFFC1111F1005FF6F1104444889D31150945F124E4B73322222225005";
constant po_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_3 ----------------------------------------------------------------------------------
constant po_3_00 : BIT_VECTOR := X"C2F0E8E840F8020B99B99999999FCCF309009209F99CEBEB06CCCCCCCCCCCCCC";
constant po_3_01 : BIT_VECTOR := X"85C988408CFFFC1E37C0189FCFCCFC20E20EF3EF66CFFCFFF33ECEF1089C0340";
constant po_3_02 : BIT_VECTOR := X"731240E64499F7400284088FFFC00E1E0189CDEF12F800EC2F8085C800EC2F80";
constant po_3_03 : BIT_VECTOR := X"5E01101FFF25F22310FCC222FF17C228D505E8C588C0EECE22F22F6C33FF37CE";
constant po_3_04 : BIT_VECTOR := X"4EEDEEC45EBEBBEE999999999B99E805E0FCD011E99E01EEEEF7CECEFFE0F211";
constant po_3_05 : BIT_VECTOR := X"37CD979F52E9D1111011DD4459FF2C9D9EEE000F4EEDEE20F4EEDEEC45EBEB0F";
constant po_3_06 : BIT_VECTOR := X"EE9EE9EE9EE9E40099999999F98008489858F188FEC899911F999090F999CD55";
constant po_3_07 : BIT_VECTOR := X"FFFFFFFFFCD999940EE9BBB088888888801F89990F12099B90B9999999999EE9";
constant po_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

end prog_mem_content;


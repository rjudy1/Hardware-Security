
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package prog_mem_content is

-- content of pe_0 ----------------------------------------------------------------------------------
constant pe_0_00 : BIT_VECTOR := X"9049A89DFA409ADEFEFFFFFFFFF88C412492595C5550AEF10840C613579BDF1F";
constant pe_0_01 : BIT_VECTOR := X"F71A99E97F333928581FF7380C06E01E31A688913210D0309001365127949FF8";
constant pe_0_02 : BIT_VECTOR := X"99C3F031F10A19E9019C318794912176FF7110690BF034F0320EF7FEB4F0320E";
constant pe_0_03 : BIT_VECTOR := X"B08D0060F64589104EB435E9B8936F58FEF700F7207220066A94D85196815101";
constant pe_0_04 : BIT_VECTOR := X"78050103F9000478FFFFFFFFDEFF27790C01004C18F00567121A68036D0F0288";
constant pe_0_05 : BIT_VECTOR := X"911A1919741FFE808AFFFF092000017805D80103F9901100178050103FB60001";
constant pe_0_06 : BIT_VECTOR := X"09D8AFFEE88D8901C40F70FD03606CF1BFF042A77AB10A7749118069306F106F";
constant pe_0_07 : BIT_VECTOR := X"2F19B950DF819BDF9BDF9C1127CFFC1B8FFDEFADFFFFFFFFF08C08F08D08608B";
constant pe_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB23";
constant pe_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_1 ----------------------------------------------------------------------------------
constant pe_1_00 : BIT_VECTOR := X"0889A8C32D8173CD0DD1FDB97426F1FEA0DA0F8003B4EDC1077768FFFFFFFF01";
constant pe_1_01 : BIT_VECTOR := X"5ABA3728F58889E29987F8F81811811011B07922211881886A1BAB8794F81424";
constant pe_1_02 : BIT_VECTOR := X"24464333868037290702970F886AA0FB3F4F09BB91F198450422391EA8450424";
constant pe_1_03 : BIT_VECTOR := X"3850B80118000E28E011A0A005A938445A5A865A86A30230A0090A821B8CA53A";
constant pe_1_04 : BIT_VECTOR := X"88980E892088C880368ACE0CCD0908FF830498EEEF0831BA0058B8901280001F";
constant pe_1_05 : BIT_VECTOR := X"0A8697A86BB976E22F008A968760928898A80E892C88D209288980E892E88092";
constant pe_1_06 : BIT_VECTOR := X"90EF80CC8118D8E0E1322239A5351282FC0A86B350970B79BA43144CB44C3323";
constant pe_1_07 : BIT_VECTOR := X"695F2BEAE0FDB1FDB9753E402AFCE85CEECCD0CCC0ECA8642908908908908908";
constant pe_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE6";
constant pe_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_2 ----------------------------------------------------------------------------------
constant pe_2_00 : BIT_VECTOR := X"411EBB17F11611FF673322222229427770770F1011103F546333333333333340";
constant pe_2_01 : BIT_VECTOR := X"F1C481F3105762E44F1AFC16864D224F04E04F0000032122040C212C0D1E0FFD";
constant pe_2_02 : BIT_VECTOR := X"4051F0EFF550E1FBC10F11016674A011AFC1001600482DF00007F1742DF00007";
constant pe_2_03 : BIT_VECTOR := X"1240E400F8000E41D0DDC0E004EDE7AEF1F101F111E0010000000EF00050EF0E";
constant pe_2_04 : BIT_VECTOR := X"8B0B0701F1080BB500000011FF6F01F02E3001DF0F13411C000D15000130004F";
constant pe_2_05 : BIT_VECTOR := X"4DDFDFDFF00FFF41010033006110008B0BF30701F001560008B0B0701F002000";
constant pe_2_06 : BIT_VECTOR := X"04E4011136711BD4107F13F1171500FD133DFF555E157555073D0DF70DF139F1";
constant pe_2_07 : BIT_VECTOR := X"0111FFF01E4D110044448F063D100951E22FF6B733222222205C057057056055";
constant pe_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB00";
constant pe_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of pe_3 ----------------------------------------------------------------------------------
constant pe_3_00 : BIT_VECTOR := X"F89288085C8800BBBB99999999969D0F1CF1929C999EEBE26CCCCCCCCCCCCCCC";
constant pe_3_01 : BIT_VECTOR := X"402280580C33380F5210EF03636F3629C29CF0CCC6633633FFE2D031EF02F452";
constant pe_3_02 : BIT_VECTOR := X"FC8D5E22499C205008C588C033F115D00EF05E00EC86D2EEC8884078D2EEC888";
constant pe_3_03 : BIT_VECTOR := X"DEFC2FCC57CCC7F80C222C7CCF22F7124040E84088FECEEC6CC6C22FFC3F22E2";
constant pe_3_04 : BIT_VECTOR := X"EBEB0F4EEDEEEBB999999999BBBEC8CDEC21E800ECDEFD0FCCF20EECCDECECFC";
constant pe_3_05 : BIT_VECTOR := X"F11011110EE44793309999EDE99C45EBEBC20F4EEDEE09C45EBEB0F4EEDEEC45";
constant pe_3_06 : BIT_VECTOR := X"E95F3990999902280C8588408088CCEF0991109992009999EF9FF52FE5209199";
constant pe_3_07 : BIT_VECTOR := X"00905CEE0B91888888888C592F099100299BBB1B999999999E9EE9EE9EE9EE9E";
constant pe_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCE0";
constant pe_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant pe_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_0 ----------------------------------------------------------------------------------
constant po_0_00 : BIT_VECTOR := X"3873F90CFE17C6CF82DFFFFFFFF0F01F3DE3D8F575570D4F0062EA92468ACE02";
constant po_0_01 : BIT_VECTOR := X"FD63A8F706911F143FFFF04121691C90A90A6A0784699C990B001011904A95F3";
constant po_0_02 : BIT_VECTOR := X"F548FEA0FF007FF7870F720791E11110FF045400803EC1F2B617FD7FC1F2B617";
constant po_0_03 : BIT_VECTOR := X"F060140039AE2EA01E4134A324BED8ACCFAE017C31870058A549A4018098F95A";
constant po_0_04 : BIT_VECTOR := X"3FA300017805010FFFFFFFFFFF82F0610693261D0AA06B0D0B16C02812064410";
constant po_0_05 : BIT_VECTOR := X"80111A8A8CEFFEF11ACF8F000320103F6209200178059E0103FC700017805010";
constant po_0_06 : BIT_VECTOR := X"8FFC18FF7C1C7192BB7F0C1F142572F34FF8539776C819776A209AF6F178E01A";
constant po_0_07 : BIT_VECTOR := X"0011FE308DEFEACE8ACE8A111048FD118BF9F8BEFFFFFFFFF8608F08708D08F0";
constant po_0_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF18";
constant po_0_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_0_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_1 ----------------------------------------------------------------------------------
constant po_1_00 : BIT_VECTOR := X"C88F99A23981F860F6CC0ECA8630F03EB1FB0EE902A1FCD18077666FFFFFFF00";
constant po_1_01 : BIT_VECTOR := X"541A4239820930F299B8688501072009EB9A1991112332653810E92868803839";
constant po_1_02 : BIT_VECTOR := X"18445A23977991398063986161EBB2094288F08BA81E5B50413F321F5B50413F";
constant po_1_03 : BIT_VECTOR := X"19B1B01AA081AAE8FFA001AA3349038514749704970F2302AA1A9A8B88718522";
constant po_1_04 : BIT_VECTOR := X"92F880928898D1882479BDF1D0F689F09B0F0BFFF4B9B49888A80908AA9BAB01";
constant po_1_05 : BIT_VECTOR := X"6297A869733A86685A8019A89660E892B880809288987C0E892D8809288980E8";
constant po_1_06 : BIT_VECTOR := X"08FF901D19091E0FF8233832B44242902D1097C240A06C68AE04444F0440D312";
constant po_1_07 : BIT_VECTOR := X"986439FB0CD0CA0ECA86425AA220D934A6D00FDDD1FDB9753089089089089089";
constant po_1_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE4";
constant po_1_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_1_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_2 ----------------------------------------------------------------------------------
constant po_2_00 : BIT_VECTOR := X"13C13B87F1F21E1E47733222222FF07372172F11D1100F0E0033333333333344";
constant po_2_01 : BIT_VECTOR := X"7F0488F1100000C00DFAA114040140FD0ED0F0DD000400404220F04CE11012F1";
constant po_2_02 : BIT_VECTOR := X"E7AEF108FF55F6F1BE1F111F50048010AA11F2246FD411F0DF017F0411F0DF01";
constant po_2_03 : BIT_VECTOR := X"F017AD7EC0DFEED3D1E00DEDCE4F0ED51F1F010F11011000EFFEDE1077046F00";
constant po_2_04 : BIT_VECTOR := X"1F0040008B0B0AFF000000011E46F510014F11DF0440140222E80007CE01ECB7";
constant po_2_05 : BIT_VECTOR := X"40DDDFFFF00FFF3117F013090000701F009430008B0B410701F0010008B0B070";
constant po_2_06 : BIT_VECTOR := X"53F1551173616655113F533F14711FF01335FF75541557555F02D30F03056D40";
constant po_2_07 : BIT_VECTOR := X"1111F1005FF6F1104444889D31150945F124E4B7332222222500560500560540";
constant po_2_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC";
constant po_2_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_2_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

-- content of po_3 ----------------------------------------------------------------------------------
constant po_3_00 : BIT_VECTOR := X"C2F0E8E840F8020B99B99999999FCCF309009209F99CEBEB06CCCCCCCCCCCCCC";
constant po_3_01 : BIT_VECTOR := X"85C988408CFFFC1E37C0189FCFCCFC20E20EF3EF66CFFCFFF33ECEF1089C0340";
constant po_3_02 : BIT_VECTOR := X"731240E64499F7400284088FFFC00E1E0189CDEF12F800EC2F8085C800EC2F80";
constant po_3_03 : BIT_VECTOR := X"5E01101FFF25F22310FCC222FF17C228D505E8C588C0EECE22F22F6C33FF37CE";
constant po_3_04 : BIT_VECTOR := X"EEDEEC45EBEBEBEE999999999B99E805E0FCD011E99E01EEEEF7CECEFFE0F211";
constant po_3_05 : BIT_VECTOR := X"9D1111011DD4459FF2C9D9EEE000F4EEDEEFBC45EBEBF30F4EEDEEC45EBEB0F4";
constant po_3_06 : BIT_VECTOR := X"9E40099999999F98008489858F188FEC899911F999090F999CD5537CD979F52E";
constant po_3_07 : BIT_VECTOR := X"999940EE9BBB088888888801F89990F12099B90B9999999999EE9EE9EE9EE9EE";
constant po_3_08 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCD";
constant po_3_09 : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0A : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0B : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0C : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0D : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0E : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
constant po_3_0F : BIT_VECTOR := X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";

end prog_mem_content;

